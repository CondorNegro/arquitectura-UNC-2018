`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Trabajo Pr�ctico N� 1. ALU.
// ALU.
// Integrantes: Kleiner Mat�as, L�pez Gast�n.
// Materia: Arquitectura de Computadoras.
// FCEFyN. UNC.
// A�o 2018.
//////////////////////////////////////////////////////////////////////////////////

// Constantes.
`define CANT_SWITCHES 6
`define CANT_BOTONES 4
`define CANT_LEDS 6

module alu(   
    i_clock,
    i_reset,  
    i_switch, 
    i_enable,
    o_leds
    );

// Par�metros.
parameter CANT_SWITCHES=`CANT_SWITCHES;
parameter CANT_BOTONES=`CANT_BOTONES;
parameter CANT_LEDS=`CANT_LEDS;

// Entradas - Salidas.
input i_clock;                              // Clock.
input [CANT_SWITCHES - 1 : 0] i_switch;     // Switches (para introducir operandos y operadores).
input i_reset;                              // Reset (hard reset).
input [CANT_BOTONES - 1 : 0] i_enable;      // Botones para indicar qu� elemento de la operaci�n es lo que se se�ala con los switches (primer operando, operador o segundo operando).
output [CANT_LEDS - 1 : 0] o_leds;          // Leds para indicar el resultado binario.

// Registros.
reg signed [CANT_SWITCHES - 1 : 0] reg_operando_1;  
reg signed [CANT_SWITCHES - 1 : 0] reg_operando_2; 
reg [CANT_SWITCHES - 1 : 0] reg_operacion;
reg signed [CANT_LEDS - 1 : 0] reg_resultado_operacion;


always@(posedge i_clock) begin
    
    //Se resetean los registros
    if (i_reset) begin
        reg_operando_1 <= 0;
        reg_operando_2 <= 0;
        reg_operacion <= 0;
        reg_resultado_operacion <= 0;
    end
    
    else begin
        //Si se presiona el boton 1 (001), se guarda el valor del switch en reg_operando_1
        if (i_enable  == 1) begin 
            reg_operando_1 <= i_switch;		
        end
        
        //Si se presiona el boton 2 (010), se guarda el valor del switch en reg_operacion.
        if (i_enable == 2) begin 
            reg_operacion <= i_switch; 	
        end
        
        //Si se presiona el boton 3 (100), se guarda el valor del switch en reg_operando_2
        if (i_enable == 4) begin  
            reg_operando_2 <= i_switch;	      
        end
        
        // De otra forma, los registros mantienen su valor.
        else begin  
            reg_operacion <= reg_operacion;
            reg_operando_1 <= reg_operando_1;	   
            reg_operando_2 <= reg_operando_2;	      
        end
    
        
        // Case donde se testea el valor de la operaci�n y en base a eso se opera entre operando1 y operando2.
        // Operaciones basadas en MIPS IV Instruction Set.
        case (reg_operacion)
            
            //ADD
            6'b100000 : begin
               reg_resultado_operacion <= reg_operando_1 + reg_operando_2;
            end
             
             //SUB
             6'b100010 : begin
               reg_resultado_operacion <= reg_operando_1 - reg_operando_2;
             end
            
            //AND
             6'b100100 : begin
                reg_resultado_operacion <= reg_operando_1 & reg_operando_2;
             end
             
             //OR
             6'b100101 : begin
                reg_resultado_operacion <= reg_operando_1 | reg_operando_2;
             end
            
            //XOR
             6'b100110 : begin
               reg_resultado_operacion <= reg_operando_1 ^ reg_operando_2;
             end
             
             //SRA (Shift Right Aritmethic).
             6'b000011 : begin
                 reg_resultado_operacion <= reg_operando_1 >>> reg_operando_2;
             end
                         
            //SRL  (Shift Right Logical).
            6'b000010 : begin
               reg_resultado_operacion <= reg_operando_1 >> reg_operando_2;
            end
            
            //NOR
            6'b100111 : begin
               reg_resultado_operacion <= ! (reg_operando_1 | reg_operando_2);
            end
            
            default : begin
                reg_resultado_operacion <= reg_resultado_operacion;
            end
            
        endcase
    end
end 

// Asignaci�n de salida.
assign {o_leds} = reg_resultado_operacion;

endmodule

