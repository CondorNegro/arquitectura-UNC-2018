`timescale 1ns / 100ps

//////////////////////////////////////////////////////////////////////////////////
// Trabajo Pr�ctico N� 1. ALU.
// Test bench de la ALU.
// Integrantes: Kleiner Mat�as, L�pez Gast�n.
// Materia: Arquitectura de Computadoras.
// FCEFyN. UNC.
// A�o 2018.
//////////////////////////////////////////////////////////////////////////////////

`define BUS_DATOS           4   // Tama�o del bus de entrada. (Por ejemplo, cantidad de switches).
`define BUS_SALIDA          4   // Tama�o del bus de salida. (Por ejemplo, cantidad de leds).
`define CANT_BOTONES_ALU    4   // Cantidad de botones.

module TestBenchAlu();
	
	
	// Par�metros
    parameter BUS_DATOS = `BUS_DATOS;
    parameter BUS_SALIDA = `BUS_SALIDA;
    parameter CANT_BOTONES_ALU = `CANT_BOTONES_ALU;
	
	//Todo puerto de salida del m�dulo es un cable.
	//Todo puerto de est�mulo o generaci�n de entrada es un registro.
	
	// Entradas - Salidas
    reg clock;                                  // Clock.
    reg hard_reset;                             // Reset.
    reg [BUS_DATOS - 1 : 0] switches;           // Switches.
    reg [CANT_BOTONES_ALU - 1 : 0] botones;     // Botones.
    wire [BUS_SALIDA - 1 : 0] leds;             // Leds.
	
	
	initial	begin
		clock = 1'b0;
		hard_reset = 1'b1; // Reset en 1.
		switches = 4'b0000; 
		botones = 4'b0000;
		#10 hard_reset = 1'b0; // Bajo el reset.
		
		// Test 1: cargar primer operando.
		#10 botones[0] = 1'b1;
		#10 switches = 4'b0101;
		#10 botones[0] = 1'b0;
		
		// Test 2: cargar segundo operando.
		#10 botones[1] = 1'b1;
        #10 switches = 4'b1000; //ADD
        #10 botones[1] = 1'b0;
		
		// Test 3: cargar tercer operando.
		#10 botones[2] = 1'b1;
        #10 switches = 4'b0101;
        #10 botones[2] = 1'b0;
		
		
		// Test 4: ADD.
		#50 botones[0] = 1'b1;
        #10 switches = 4'b1101;
        #10 botones[0] = 1'b0;
        #10 botones[1] = 1'b1;
        #10 switches = 4'b1000; //ADD
        #10 botones[1] = 1'b0;
        #10 botones[2] = 1'b1;
        #10 switches = 4'b0101;
        #10 botones[2] = 1'b0;
		
		
		// Test 5: SUB.
		#50 botones[0] = 1'b1;
        #10 switches = 4'b0101;
        #10 botones[0] = 1'b0;
        #10 botones[1] = 1'b1;
        #10 switches = 4'b1010; //SUB
        #10 botones[1] = 1'b0;
        #10 botones[2] = 1'b1;
        #10 switches = 4'b0001;
        #10 botones[2] = 1'b0;
		
		
		// Test 6: AND.
        #50 botones[0] = 1'b1;
        #10 switches = 4'b1101;
        #10 botones[0] = 1'b0;
        #10 botones[1] = 1'b1;
        #10 switches = 4'b1100; //AND
        #10 botones[1] = 1'b0;
        #10 botones[2] = 1'b1;
        #10 switches = 4'b0101;
        #10 botones[2] = 1'b0;        
        
        
        // Test 7: OR.
         #50 botones[0] = 1'b1;
         #10 switches = 4'b1101;
         #10 botones[0] = 1'b0;
         #10 botones[1] = 1'b1;
         #10 switches = 4'b1101; //OR
         #10 botones[1] = 1'b0;
         #10 botones[2] = 1'b1;
         #10 switches = 4'b0101;
         #10 botones[2] = 1'b0;       
		
        // Test 8: XOR.
         #50 botones[0] = 1'b1;
         #10 switches = 4'b1101;
         #10 botones[0] = 1'b0;
         #10 botones[1] = 1'b1;
         #10 switches = 4'b1110; //XOR
         #10 botones[1] = 1'b0;
         #10 botones[2] = 1'b1;
         #10 switches = 4'b0101;
         #10 botones[2] = 1'b0;       
          
                
        // Test 9: SRA.
		 #50 botones[0] = 1'b1;
         #10 switches = 4'b1101;
         #10 botones[0] = 1'b0;
         #10 botones[1] = 1'b1;
         #10 switches = 4'b0011; //SRA
         #10 botones[1] = 1'b0;
         #10 botones[2] = 1'b1;
         #10 switches = 4'b0011;
         #10 botones[2] = 1'b0;       
		
		// Test 10: SRL.
		 #50 botones[0] = 1'b1;
         #10 switches = 4'b1101;
         #10 botones[0] = 1'b0;
         #10 botones[1] = 1'b1;
         #10 switches = 4'b0010; //SRL
         #10 botones[1] = 1'b0;
         #10 botones[2] = 1'b1;
         #10 switches = 4'b0011;
         #10 botones[2] = 1'b0;       
		
		// Test 11: NOR.
		 #50 botones[0] = 1'b1;
         #10 switches = 4'b1101;
         #10 botones[0] = 1'b0;
         #10 botones[1] = 1'b1;
         #10 switches = 4'b1111; //NOR
         #10 botones[1] = 1'b0;
         #10 botones[2] = 1'b1;
         #10 switches = 4'b0101;
         #10 botones[2] = 1'b0;       
		
		// Test 12: Operaci�n falsa.
        #50 botones[0] = 1'b1;
        #10 switches = 4'b1101;
        #10 botones[0] = 1'b0;
        #10 botones[1] = 1'b1;
        #10 switches = 4'b0000; //Falsa.
        #10 botones[1] = 1'b0;
        #10 botones[2] = 1'b1;
        #10 switches = 4'b0101;
        #10 botones[2] = 1'b0;      
		
		// Test 13: Prueba reset.
		#100 hard_reset = 1'b1; // Reset.
		#10 hard_reset = 1'b0; // Bajo el reset.
		
		
		#1000000000 $finish;
	end
	
	always #2.5 clock=~clock;  // Simulaci�n de clock.



//M�dulo para pasarle los est�mulos del banco de pruebas.
alu
    #(
         .CANT_SWITCHES (BUS_DATOS),
         .CANT_LEDS (BUS_SALIDA),
         .CANT_BOTONES (CANT_BOTONES_ALU)
     ) 
   u_alu1    // Una sola instancia de este m�dulo
   (
   .i_clock (clock),
   .i_reset (hard_reset),
   .i_switch (switches),
   .i_enable (botones),
   .o_leds (leds)
   );
   
endmodule

